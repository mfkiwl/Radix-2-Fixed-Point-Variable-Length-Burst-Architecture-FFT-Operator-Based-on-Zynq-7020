`timescale 1ns / 1ps

module tb_fft_top_new;

  // Parameters
  parameter CLK_PERIOD = 10;  // Clock period in ns (100 MHz)

  // Testbench signals
  reg         i_clk;
  reg         i_rst_n;
  reg         i_n_cfg_valid;
  reg  [4:0]  i_n_cfg;
  reg         i_data_in_valid;
  reg  [31:0] i_data_in;

  wire [31:0] o_data_out;
  wire        o_data_out_valid;
  wire        o_idle_out;
  reg [5:0] n;


  // Instantiate the fft_top module
  fft_top_new uut (
                .i_clk(i_clk),
                .i_rst_n(i_rst_n),
                .i_n_cfg_valid(i_n_cfg_valid),
                .i_n_cfg(i_n_cfg),
                .i_data_in_valid(i_data_in_valid),
                .i_data_in(i_data_in),
                .o_data_out(o_data_out),
                .o_data_out_valid(o_data_out_valid),
                .o_idle_out(o_idle_out)
              );

  integer i;
  integer output_file;
  reg [8*255:0] filename;

  // Clock generation
  initial
  begin
    i_clk = 0;
    forever
      #(CLK_PERIOD / 2) i_clk = ~i_clk;
  end

  /*
    //debugging ports
    reg [15:0] i_data_in_real;
    reg [15:0] i_data_in_imag;
    always @ (posedge i_clk)
    begin
      i_data_in_real = i_data_in[31:16];
      i_data_in_imag = i_data_in[15:0];
    end
  */


  // FFT Test Configuration
  // Sample Frequency (f): 10000000 Hz
  // Phase (phi): 0.0 rad
  // Number of Samples (num_samples): 8
  // Task to configure FFT and send data
  task fft_sintest8(
      input [4:0] n_cfg        // FFT configuration value
    );
    begin
      // Start FFT configuration
      
      
      

      // Wait before sending data
      //#20;
      // Start sending data

      @(posedge i_clk);
      i_n_cfg_valid = 1;
      i_n_cfg = n_cfg;
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1

      @(posedge i_clk);
      i_n_cfg_valid = 0;
      i_n_cfg = 5'd0;
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 2

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 3

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 4

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 5

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 6

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 7

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 8

      // Stop sending data
      @(posedge i_clk);
      i_data_in_valid = 0;
      i_data_in = 32'd0;
      #(800);
    end
  endtask


  // FFT Test Configuration
  // Sample Frequency (f): 10000000 Hz
  // Phase (phi): 0.0 rad
  // Number of Samples (num_samples): 128

  // Task to configure FFT and send data
  task fft_sintest128(
      input [4:0] n_cfg        // FFT configuration value
    );
    begin
      // Start FFT configuration
      i_n_cfg_valid = 1;
      i_n_cfg = n_cfg;
      #10;
      i_n_cfg_valid = 0;
      i_n_cfg = 5'd0;

      // Wait before sending data
      #20;
      // Start sending data

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 2

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 3

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 4

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 5

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 6

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 7

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 8

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 9

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 10

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 11

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 12

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 13

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 14

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 15

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 16

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 17

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 18

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 19

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 20

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 21

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 22

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 23

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 24

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 25

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 26

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 27

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 28

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 29

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 30

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 31

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 32

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 33

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 34

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 35

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 36

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 37

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 38

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 39

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 40

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 41

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 42

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 43

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 44

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 45

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 46

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 47

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 48

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 49

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 50

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 51

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 52

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 53

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 54

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 55

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 56

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 57

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 58

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 59

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 60

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 61

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 62

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 63

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 64

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 65

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 66

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 67

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 68

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 69

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 70

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 71

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 72

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 73

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 74

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 75

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 76

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 77

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 78

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 79

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 80

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 81

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 82

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 83

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 84

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 85

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 86

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 87

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 88

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 89

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 90

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 91

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 92

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 93

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 94

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 95

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 96

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 97

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 98

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 99

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 100

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 101

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 102

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 103

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 104

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 105

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 106

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 107

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 108

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 109

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 110

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 111

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 112

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 113

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 114

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 115

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 116

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 117

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 118

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 119

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 120

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 121

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 122

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 123

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 124

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 125

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 126

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 127

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 128

      // Stop sending data
      @(posedge i_clk);
      i_data_in_valid = 0;
      i_data_in = 32'd0;
      #(8000);
    end
  endtask



  // FFT Test Configuration
  // Sample Frequency (f): 10000000 Hz
  // Phase (phi): 0.0 rad
  // Number of Samples (num_samples): 2048

  // Task to configure FFT and send data
  task fft_sintest2048(
      input [4:0] n_cfg        // FFT configuration value
    );
    begin
      // Start FFT configuration
      i_n_cfg_valid = 1;
      i_n_cfg = n_cfg;
      #10;
      i_n_cfg_valid = 0;
      i_n_cfg = 5'd0;

      // Wait before sending data
      #20;
      // Start sending data

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 2

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 3

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 4

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 5

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 6

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 7

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 8

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 9

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 10

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 11

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 12

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 13

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 14

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 15

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 16

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 17

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 18

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 19

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 20

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 21

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 22

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 23

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 24

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 25

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 26

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 27

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 28

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 29

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 30

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 31

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 32

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 33

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 34

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 35

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 36

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 37

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 38

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 39

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 40

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 41

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 42

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 43

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 44

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 45

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 46

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 47

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 48

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 49

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 50

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 51

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 52

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 53

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 54

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 55

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 56

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 57

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 58

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 59

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 60

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 61

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 62

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 63

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 64

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 65

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 66

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 67

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 68

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 69

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 70

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 71

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 72

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 73

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 74

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 75

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 76

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 77

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 78

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 79

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 80

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 81

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 82

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 83

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 84

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 85

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 86

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 87

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 88

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 89

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 90

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 91

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 92

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 93

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 94

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 95

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 96

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 97

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 98

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 99

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 100

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 101

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 102

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 103

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 104

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 105

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 106

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 107

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 108

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 109

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 110

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 111

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 112

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 113

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 114

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 115

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 116

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 117

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 118

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 119

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 120

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 121

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 122

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 123

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 124

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 125

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 126

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 127

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 128

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 129

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 130

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 131

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 132

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 133

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 134

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 135

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 136

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 137

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 138

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 139

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 140

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 141

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 142

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 143

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 144

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 145

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 146

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 147

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 148

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 149

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 150

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 151

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 152

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 153

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 154

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 155

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 156

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 157

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 158

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 159

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 160

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 161

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 162

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 163

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 164

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 165

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 166

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 167

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 168

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 169

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 170

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 171

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 172

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 173

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 174

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 175

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 176

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 177

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 178

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 179

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 180

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 181

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 182

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 183

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 184

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 185

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 186

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 187

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 188

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 189

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 190

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 191

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 192

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 193

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 194

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 195

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 196

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 197

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 198

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 199

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 200

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 201

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 202

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 203

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 204

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 205

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 206

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 207

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 208

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 209

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 210

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 211

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 212

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 213

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 214

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 215

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 216

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 217

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 218

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 219

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 220

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 221

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 222

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 223

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 224

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 225

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 226

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 227

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 228

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 229

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 230

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 231

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 232

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 233

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 234

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 235

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 236

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 237

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 238

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 239

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 240

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 241

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 242

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 243

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 244

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 245

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 246

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 247

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 248

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 249

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 250

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 251

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 252

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 253

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 254

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 255

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 256

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 257

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 258

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 259

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 260

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 261

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 262

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 263

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 264

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 265

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 266

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 267

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 268

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 269

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 270

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 271

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 272

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 273

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 274

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 275

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 276

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 277

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 278

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 279

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 280

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 281

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 282

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 283

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 284

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 285

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 286

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 287

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 288

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 289

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 290

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 291

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 292

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 293

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 294

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 295

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 296

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 297

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 298

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 299

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 300

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 301

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 302

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 303

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 304

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 305

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 306

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 307

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 308

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 309

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 310

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 311

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 312

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 313

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 314

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 315

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 316

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 317

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 318

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 319

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 320

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 321

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 322

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 323

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 324

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 325

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 326

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 327

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 328

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 329

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 330

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 331

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 332

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 333

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 334

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 335

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 336

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 337

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 338

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 339

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 340

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 341

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 342

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 343

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 344

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 345

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 346

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 347

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 348

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 349

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 350

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 351

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 352

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 353

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 354

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 355

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 356

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 357

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 358

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 359

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 360

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 361

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 362

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 363

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 364

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 365

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 366

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 367

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 368

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 369

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 370

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 371

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 372

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 373

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 374

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 375

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 376

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 377

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 378

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 379

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 380

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 381

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 382

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 383

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 384

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 385

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 386

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 387

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 388

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 389

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 390

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 391

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 392

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 393

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 394

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 395

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 396

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 397

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 398

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 399

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 400

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 401

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 402

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 403

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 404

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 405

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 406

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 407

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 408

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 409

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 410

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 411

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 412

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 413

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 414

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 415

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 416

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 417

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 418

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 419

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 420

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 421

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 422

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 423

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 424

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 425

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 426

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 427

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 428

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 429

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 430

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 431

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 432

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 433

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 434

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 435

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 436

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 437

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 438

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 439

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 440

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 441

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 442

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 443

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 444

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 445

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 446

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 447

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 448

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 449

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 450

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 451

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 452

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 453

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 454

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 455

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 456

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 457

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 458

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 459

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 460

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 461

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 462

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 463

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 464

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 465

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 466

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 467

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 468

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 469

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 470

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 471

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 472

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 473

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 474

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 475

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 476

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 477

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 478

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 479

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 480

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 481

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 482

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 483

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 484

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 485

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 486

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 487

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 488

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 489

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 490

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 491

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 492

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 493

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 494

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 495

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 496

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 497

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 498

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 499

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 500

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 501

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 502

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 503

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 504

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 505

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 506

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 507

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 508

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 509

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 510

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 511

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 512

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 513

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 514

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 515

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 516

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 517

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 518

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 519

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 520

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 521

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 522

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 523

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 524

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 525

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 526

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 527

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 528

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 529

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 530

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 531

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 532

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 533

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 534

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 535

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 536

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 537

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 538

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 539

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 540

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 541

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 542

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 543

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 544

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 545

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 546

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 547

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 548

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 549

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 550

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 551

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 552

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 553

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 554

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 555

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 556

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 557

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 558

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 559

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 560

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 561

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 562

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 563

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 564

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 565

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 566

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 567

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 568

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 569

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 570

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 571

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 572

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 573

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 574

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 575

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 576

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 577

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 578

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 579

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 580

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 581

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 582

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 583

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 584

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 585

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 586

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 587

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 588

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 589

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 590

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 591

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 592

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 593

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 594

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 595

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 596

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 597

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 598

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 599

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 600

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 601

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 602

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 603

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 604

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 605

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 606

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 607

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 608

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 609

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 610

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 611

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 612

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 613

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 614

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 615

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 616

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 617

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 618

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 619

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 620

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 621

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 622

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 623

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 624

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 625

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 626

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 627

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 628

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 629

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 630

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 631

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 632

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 633

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 634

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 635

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 636

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 637

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 638

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 639

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 640

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 641

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 642

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 643

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 644

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 645

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 646

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 647

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 648

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 649

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 650

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 651

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 652

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 653

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 654

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 655

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 656

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 657

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 658

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 659

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 660

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 661

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 662

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 663

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 664

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 665

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 666

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 667

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 668

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 669

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 670

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 671

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 672

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 673

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 674

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 675

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 676

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 677

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 678

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 679

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 680

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 681

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 682

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 683

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 684

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 685

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 686

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 687

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 688

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 689

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 690

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 691

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 692

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 693

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 694

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 695

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 696

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 697

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 698

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 699

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 700

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 701

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 702

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 703

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 704

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 705

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 706

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 707

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 708

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 709

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 710

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 711

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 712

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 713

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 714

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 715

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 716

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 717

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 718

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 719

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 720

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 721

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 722

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 723

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 724

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 725

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 726

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 727

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 728

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 729

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 730

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 731

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 732

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 733

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 734

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 735

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 736

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 737

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 738

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 739

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 740

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 741

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 742

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 743

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 744

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 745

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 746

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 747

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 748

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 749

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 750

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 751

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 752

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 753

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 754

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 755

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 756

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 757

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 758

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 759

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 760

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 761

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 762

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 763

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 764

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 765

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 766

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 767

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 768

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 769

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 770

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 771

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 772

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 773

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 774

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 775

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 776

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 777

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 778

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 779

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 780

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 781

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 782

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 783

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 784

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 785

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 786

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 787

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 788

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 789

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 790

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 791

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 792

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 793

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 794

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 795

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 796

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 797

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 798

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 799

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 800

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 801

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 802

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 803

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 804

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 805

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 806

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 807

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 808

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 809

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 810

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 811

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 812

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 813

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 814

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 815

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 816

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 817

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 818

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 819

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 820

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 821

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 822

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 823

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 824

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 825

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 826

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 827

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 828

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 829

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 830

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 831

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 832

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 833

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 834

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 835

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 836

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 837

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 838

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 839

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 840

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 841

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 842

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 843

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 844

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 845

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 846

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 847

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 848

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 849

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 850

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 851

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 852

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 853

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 854

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 855

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 856

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 857

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 858

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 859

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 860

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 861

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 862

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 863

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 864

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 865

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 866

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 867

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 868

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 869

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 870

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 871

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 872

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 873

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 874

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 875

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 876

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 877

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 878

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 879

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 880

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 881

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 882

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 883

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 884

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 885

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 886

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 887

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 888

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 889

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 890

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 891

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 892

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 893

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 894

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 895

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 896

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 897

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 898

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 899

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 900

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 901

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 902

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 903

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 904

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 905

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 906

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 907

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 908

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 909

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 910

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 911

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 912

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 913

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 914

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 915

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 916

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 917

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 918

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 919

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 920

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 921

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 922

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 923

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 924

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 925

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 926

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 927

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 928

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 929

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 930

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 931

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 932

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 933

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 934

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 935

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 936

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 937

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 938

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 939

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 940

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 941

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 942

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 943

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 944

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 945

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 946

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 947

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 948

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 949

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 950

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 951

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 952

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 953

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 954

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 955

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 956

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 957

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 958

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 959

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 960

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 961

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 962

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 963

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 964

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 965

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 966

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 967

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 968

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 969

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 970

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 971

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 972

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 973

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 974

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 975

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 976

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 977

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 978

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 979

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 980

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 981

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 982

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 983

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 984

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 985

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 986

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 987

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 988

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 989

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 990

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 991

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 992

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 993

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 994

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 995

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 996

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 997

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 998

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 999

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1000

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1001

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1002

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1003

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1004

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1005

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1006

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1007

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1008

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1009

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1010

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1011

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1012

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1013

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1014

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1015

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1016

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1017

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1018

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1019

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1020

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1021

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1022

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1023

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1024

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1025

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1026

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1027

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1028

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1029

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1030

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1031

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1032

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1033

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1034

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1035

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1036

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1037

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1038

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1039

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1040

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1041

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1042

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1043

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1044

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1045

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1046

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1047

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1048

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1049

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1050

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1051

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1052

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1053

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1054

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1055

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1056

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1057

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1058

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1059

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1060

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1061

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1062

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1063

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1064

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1065

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1066

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1067

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1068

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1069

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1070

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1071

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1072

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1073

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1074

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1075

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1076

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1077

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1078

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1079

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1080

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1081

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1082

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1083

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1084

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1085

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1086

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1087

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1088

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1089

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1090

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1091

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1092

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1093

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1094

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1095

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1096

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1097

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1098

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1099

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1100

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1101

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1102

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1103

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1104

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1105

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1106

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1107

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1108

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1109

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1110

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1111

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1112

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1113

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1114

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1115

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1116

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1117

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1118

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1119

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1120

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1121

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1122

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1123

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1124

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1125

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1126

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1127

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1128

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1129

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1130

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1131

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1132

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1133

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1134

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1135

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1136

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1137

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1138

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1139

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1140

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1141

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1142

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1143

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1144

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1145

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1146

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1147

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1148

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1149

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1150

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1151

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1152

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1153

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1154

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1155

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1156

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1157

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1158

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1159

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1160

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1161

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1162

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1163

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1164

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1165

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1166

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1167

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1168

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1169

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1170

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1171

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1172

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1173

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1174

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1175

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1176

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1177

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1178

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1179

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1180

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1181

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1182

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1183

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1184

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1185

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1186

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1187

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1188

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1189

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1190

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1191

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1192

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1193

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1194

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1195

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1196

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1197

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1198

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1199

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1200

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1201

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1202

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1203

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1204

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1205

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1206

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1207

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1208

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1209

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1210

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1211

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1212

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1213

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1214

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1215

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1216

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1217

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1218

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1219

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1220

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1221

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1222

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1223

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1224

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1225

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1226

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1227

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1228

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1229

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1230

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1231

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1232

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1233

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1234

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1235

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1236

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1237

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1238

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1239

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1240

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1241

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1242

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1243

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1244

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1245

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1246

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1247

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1248

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1249

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1250

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1251

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1252

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1253

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1254

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1255

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1256

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1257

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1258

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1259

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1260

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1261

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1262

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1263

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1264

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1265

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1266

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1267

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1268

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1269

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1270

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1271

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1272

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1273

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1274

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1275

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1276

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1277

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1278

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1279

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1280

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1281

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1282

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1283

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1284

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1285

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1286

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1287

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1288

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1289

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1290

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1291

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1292

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1293

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1294

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1295

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1296

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1297

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1298

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1299

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1300

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1301

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1302

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1303

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1304

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1305

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1306

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1307

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1308

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1309

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1310

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1311

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1312

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1313

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1314

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1315

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1316

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1317

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1318

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1319

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1320

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1321

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1322

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1323

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1324

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1325

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1326

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1327

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1328

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1329

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1330

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1331

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1332

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1333

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1334

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1335

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1336

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1337

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1338

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1339

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1340

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1341

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1342

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1343

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1344

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1345

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1346

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1347

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1348

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1349

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1350

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1351

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1352

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1353

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1354

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1355

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1356

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1357

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1358

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1359

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1360

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1361

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1362

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1363

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1364

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1365

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1366

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1367

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1368

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1369

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1370

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1371

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1372

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1373

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1374

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1375

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1376

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1377

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1378

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1379

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1380

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1381

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1382

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1383

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1384

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1385

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1386

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1387

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1388

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1389

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1390

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1391

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1392

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1393

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1394

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1395

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1396

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1397

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1398

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1399

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1400

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1401

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1402

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1403

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1404

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1405

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1406

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1407

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1408

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1409

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1410

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1411

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1412

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1413

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1414

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1415

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1416

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1417

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1418

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1419

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1420

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1421

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1422

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1423

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1424

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1425

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1426

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1427

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1428

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1429

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1430

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1431

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1432

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1433

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1434

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1435

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1436

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1437

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1438

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1439

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1440

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1441

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1442

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1443

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1444

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1445

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1446

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1447

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1448

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1449

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1450

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1451

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1452

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1453

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1454

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1455

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1456

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1457

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1458

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1459

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1460

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1461

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1462

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1463

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1464

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1465

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1466

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1467

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1468

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1469

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1470

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1471

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1472

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1473

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1474

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1475

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1476

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1477

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1478

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1479

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1480

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1481

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1482

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1483

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1484

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1485

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1486

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1487

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1488

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1489

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1490

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1491

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1492

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1493

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1494

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1495

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1496

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1497

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1498

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1499

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1500

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1501

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1502

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1503

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1504

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1505

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1506

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1507

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1508

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1509

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1510

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1511

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1512

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1513

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1514

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1515

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1516

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1517

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1518

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1519

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1520

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1521

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1522

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1523

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1524

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1525

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1526

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1527

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1528

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1529

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1530

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1531

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1532

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1533

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1534

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1535

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1536

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1537

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1538

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1539

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1540

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1541

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1542

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1543

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1544

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1545

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1546

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1547

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1548

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1549

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1550

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1551

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1552

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1553

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1554

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1555

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1556

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1557

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1558

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1559

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1560

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1561

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1562

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1563

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1564

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1565

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1566

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1567

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1568

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1569

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1570

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1571

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1572

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1573

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1574

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1575

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1576

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1577

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1578

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1579

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1580

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1581

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1582

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1583

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1584

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1585

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1586

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1587

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1588

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1589

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1590

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1591

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1592

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1593

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1594

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1595

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1596

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1597

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1598

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1599

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1600

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1601

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1602

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1603

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1604

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1605

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1606

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1607

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1608

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1609

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1610

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1611

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1612

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1613

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1614

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1615

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1616

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1617

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1618

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1619

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1620

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1621

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1622

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1623

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1624

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1625

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1626

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1627

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1628

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1629

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1630

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1631

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1632

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1633

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1634

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1635

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1636

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1637

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1638

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1639

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1640

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1641

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1642

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1643

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1644

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1645

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1646

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1647

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1648

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1649

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1650

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1651

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1652

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1653

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1654

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1655

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1656

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1657

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1658

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1659

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1660

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1661

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1662

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1663

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1664

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1665

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1666

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1667

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1668

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1669

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1670

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1671

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1672

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1673

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1674

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1675

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1676

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1677

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1678

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1679

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1680

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1681

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1682

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1683

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1684

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1685

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1686

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1687

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1688

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1689

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1690

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1691

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1692

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1693

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1694

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1695

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1696

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1697

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1698

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1699

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1700

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1701

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1702

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1703

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1704

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1705

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1706

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1707

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1708

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1709

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1710

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1711

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1712

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1713

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1714

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1715

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1716

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1717

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1718

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1719

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1720

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1721

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1722

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1723

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1724

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1725

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1726

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1727

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1728

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1729

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1730

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1731

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1732

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1733

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1734

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1735

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1736

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1737

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1738

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1739

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1740

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1741

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1742

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1743

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1744

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1745

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1746

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1747

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1748

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1749

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1750

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1751

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1752

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1753

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1754

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1755

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1756

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1757

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1758

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1759

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1760

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1761

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1762

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1763

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1764

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1765

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1766

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1767

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1768

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1769

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1770

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1771

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1772

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1773

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1774

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1775

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1776

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1777

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1778

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1779

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1780

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1781

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1782

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1783

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1784

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1785

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1786

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1787

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1788

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1789

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1790

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1791

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1792

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1793

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1794

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1795

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1796

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1797

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1798

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1799

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1800

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1801

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1802

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1803

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1804

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1805

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1806

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1807

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1808

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1809

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1810

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1811

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1812

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1813

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1814

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1815

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1816

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1817

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1818

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1819

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1820

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1821

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1822

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1823

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1824

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1825

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1826

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1827

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1828

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1829

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1830

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1831

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1832

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1833

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1834

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1835

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1836

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1837

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1838

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1839

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1840

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1841

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1842

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1843

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1844

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1845

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1846

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1847

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1848

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1849

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1850

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1851

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1852

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1853

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1854

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1855

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1856

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1857

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1858

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1859

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1860

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1861

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1862

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1863

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1864

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1865

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1866

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1867

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1868

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1869

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1870

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1871

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1872

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1873

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1874

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1875

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1876

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1877

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1878

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1879

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1880

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1881

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1882

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1883

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1884

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1885

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1886

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1887

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1888

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1889

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1890

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1891

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1892

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1893

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1894

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1895

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1896

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1897

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1898

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1899

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1900

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1901

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1902

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1903

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1904

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1905

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1906

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1907

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1908

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1909

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1910

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1911

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1912

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1913

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1914

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1915

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1916

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1917

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1918

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1919

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1920

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1921

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1922

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1923

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1924

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1925

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1926

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1927

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1928

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1929

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1930

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1931

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1932

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1933

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1934

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1935

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1936

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1937

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1938

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1939

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1940

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1941

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1942

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1943

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1944

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1945

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1946

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1947

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1948

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1949

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1950

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1951

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1952

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1953

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1954

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1955

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1956

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1957

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1958

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1959

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1960

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1961

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1962

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1963

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1964

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1965

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1966

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1967

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1968

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1969

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1970

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1971

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1972

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1973

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1974

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1975

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1976

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1977

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1978

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1979

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1980

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1981

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1982

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1983

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1984

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1985

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1986

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1987

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1988

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1989

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 1990

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 1991

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 1992

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 1993

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 1994

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 1995

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 1996

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 1997

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 1998

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 1999

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 2000

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 2001

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 2002

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 2003

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 2004

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 2005

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 2006

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 2007

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 2008

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 2009

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 2010

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 2011

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 2012

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 2013

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 2014

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 2015

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 2016

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 2017

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 2018

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 2019

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 2020

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 2021

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 2022

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 2023

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 2024

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 2025

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 2026

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 2027

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 2028

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 2029

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 2030

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 2031

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 2032

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 2033

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 2034

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 2035

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 2036

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 2037

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 2038

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b1000011001000100};  // sample 2039

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b1011010011000011};  // sample 2040

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0111111111111111, 16'b0000000000000000};  // sample 2041

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0110011110001110, 16'b0100101100111101};  // sample 2042

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b0010011110001110, 16'b0111100110111100};  // sample 2043

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b0111100110111100};  // sample 2044

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b0100101100111101};  // sample 2045

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1000000000000000, 16'b0000000000000000};  // sample 2046

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1001100001110010, 16'b1011010011000011};  // sample 2047

      @(posedge i_clk);
      i_data_in_valid = 1;
      i_data_in = {16'b1101100001110010, 16'b1000011001000100};  // sample 2048

      // Stop sending data
      @(posedge i_clk);
      i_data_in_valid = 0;
      i_data_in = 32'd0;
      #(400000);
    end
  endtask



  initial
  begin
    // Initialize inputs
    i_rst_n = 0;
    i_n_cfg_valid = 0;
    i_n_cfg = 5'd0;
    i_data_in_valid = 0;
    i_data_in = 32'd0;
    // Apply reset
    #20;
    i_rst_n = 1;
    // Wait for some time after reset
    #20;

    //round1,8点
    // 定义输出文件名称
    filename = {"D:/fpga/fft_top_new/results/hw_fft_output8", ".txt"};
    // Open the output file for writing
    output_file = $fopen(filename, "wb");
    // Execute FFT test
    n = 5'd3;
    fft_sintest8(n);
    // Close the file
    $fclose(output_file);
    $finish;


    

    //round2,128点
    // 定义输出文件名称
    filename = {"D:/fpga/fft_top_new/results/hw_fft_output128", ".txt"};
    // Open the output file for writing
    output_file = $fopen(filename, "wb");
    n= 5'd7;
    // Execute FFT test
    fft_sintest128(n);
    // Close the file
    $fclose(output_file);

    //round3,2048点
    // 定义输出文件名称
    filename = {"D:/fpga/fft_top_new/results/hw_fft_output2048", ".txt"};
    // Open the output file for writing
    output_file = $fopen(filename, "wb");
    n= 5'd11;
    // Execute FFT test
    fft_sintest2048(n);
    // Close the file
    $fclose(output_file);
    



  end

  // Declare real and imaginary parts for writing binary data to file

  reg signed [15:0] real_part;
  reg signed [15:0] imag_part;


  // Monitor outputs and write to file when o_data_out_valid = 1
  always @(posedge i_clk)
  begin
    if (o_data_out_valid)
    begin
      // Extract real and imaginary parts
      real_part = o_data_out[31:16];  // Extract real part (upper 16 bits)
      imag_part = o_data_out[15:0];   // Extract imaginary part (lower 16 bits)

      // Write to file as binary with labels for real and imag
      // Write real part
      $fwrite(output_file, "%b ", real_part);
      // Write imaginary part
      $fwrite(output_file, "%b\n", imag_part);

      // Convert to decimal using q3_12_to_real function and display
      $display("Real Part (decimal): %f", q3_12_to_real(real_part));
      $display("Imaginary Part (decimal): %f", q3_12_to_real(imag_part));
    end
  end

  // Task: Convert Q3.12 format value to decimal
  function real q3_12_to_real;
    input signed [15:0] value;
    begin
      q3_12_to_real = value / 4096.0; // 2^12 = 4096
    end
  endfunction



endmodule
